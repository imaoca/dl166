 module ram(clk, we, r_addr, r_data, w_addr, w_data); 
             input clk, we;
             input  [7:0] r_addr, w_addr;
             input  [7:0] w_data;
             output [7:0] r_data;
             reg [7:0] mem [255:0];     
	     initial begin
		　mem[0] <= 8'b01100_000;// inc R0
		　mem[1] <= 8'b1000_0000;// jnc 0
		　mem[2] <= 8'b1010_0000;// MVI 0
		　mem[3] <= 8'b1001_0000;// jmp 0
	     end
             always @(posedge clk) begin
                 if(we) mem[w_addr] <= w_data; 
             end
             assign r_data = mem[r_addr];
 endmodule
